`timescale 1ns / 1ps

module ROM (
    input  logic [31:0] addr,
    output logic [31:0] data
);
    logic [31:0] rom[0:2**8-1];

    initial begin
        $readmemh("/home/aedu46/AI_HW_Verilog/RV32I_Project/TB/code.mem", rom);
    end

    // initial begin
    // //rom[x]=32'b fucn7 _ rs2 _ rs1 _f3 _ rd  _ op // R-Type
    // // rom[0] = 32'b0000000_00001_00010_000_00100_0110011;// add x4, x2, x1 O
    // // rom[1] = 32'b0100000_00001_00010_000_00101_0110011;// sub x5, x2, x1 O
    // //rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ op // I-Type
    // rom[0] = 32'h4080d213;// srai x4, x1, 8
    // rom[1] = 32'h0080d293;// srli x5, x1, 8
    // rom[2] = 32'b0000000_00000_00001_010_00110_0110011;// slt   x6, x1, x0 
    // rom[3] = 32'b0000000_00000_00001_011_00111_0110011;// sltu  x7, x1, x0
    // //rom[x]=32'b imm7  _ rs2 _ rs1 _f3 _ imm5_ op // S-Type
    // // rom[3] = 32'b0000000_00011_00000_010_01000_0100011;// sw x3, 8(x0)
    // //rom[x]=32'b imm7  _ rs2 _ rs1 _f3 _ imm5_ op // S-Type
    // rom[4] = 32'b0000000_11111_00000_010_00000_0100011;// sw x31, 0(x0)
    // //rom[x]=32'b imm[20][10:1][11][19:12]      _ rd  _ op // J-Type
    // // rom[4] = 32'b0_0000000110_0_00000000_00001_1101111;// jal x1, 12
    // //rom[x]=32'b imm[11:0]_rs1 _000_ rd  _ op // JL-Type
    // // rom[4] = 32'b000000010000_00010_000_00001_1100111;// jalr x1, x2, 16
    // //rom[x]=32'b imm7  _ rs2 _ rs1 _f3 _ imm5_ op // B-Type
    // rom[5] = 32'h0001e663;// bltu x3, x0, 12
    // // rom[6] = 32'h0001c663;// blt x3, x0, 12
    // //rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ op // L-Type
    // rom[6] = 32'b000000000000_00000_010_10111_0000011;// lw x23, 0(x0)   
    // //rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ op // I-Type
    // rom[7] = 32'b000000000001_00001_000_01001_0010011;// addi x9, x1, 1 
    // // rom[7] = 32'b000000001100_00010_000_00001_1100111;// jalr x1, x2, 12
    // rom[8] = 32'b000000000100_00010_111_01010_0010011;// andi x10, x2, 4 
    // rom[9] = 32'b000000000001_00010_110_01011_0010011;// ori x11, x2, 1 
    // // rom[10] = 32'b000000000011_00001_001_01100_0010011;// slli x12, x1, 1 // 2b00001011 << 3
    // //rom[x]=32'b imm20      _ rd  _ op // LU-Type
    // rom[10] = 32'b10000000000000000000_00101_0110111;// lui x5, 0x10000
    // //rom[x]=32'b imm20      _ rd  _ op // AU-Type
    // rom[11] = 32'b10000000000000000000_00101_0010111;// auipc x5, 0x10000
    // //rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ op // L-Type
    // rom[12] = 32'b000000000000_00000_000_01111_0000011;// lb x15, 0(x0)
    // rom[13] = 32'b000000000001_00000_000_10000_0000011;// lb x16, 1(x0)
    // rom[14] = 32'b000000000010_00000_000_10001_0000011;// lb x17, 2(x0)
    // rom[15] = 32'b000000000011_00000_000_10010_0000011;// lb x18, 3(x0)
    // //rom[x]=32'b imm7  _ rs2 _ rs1 _f3 _ imm5_ op // S-Type
    // rom[16] = 32'b0000000_11111_00001_000_00000_0100011;// sb x31, 0(x1)
    // rom[17] = 32'b0000000_11111_00001_000_00001_0100011;// sb x31, 1(x1)
    // rom[18] = 32'b0000000_11111_00001_000_00010_0100011;// sb x31, 2(x1)
    // rom[19] = 32'b0000000_11111_00001_000_00011_0100011;// sb x31, 3(x1)
    // //rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ op // L-Type
    // rom[20] = 32'b000000000000_00000_001_10011_0000011;// lh x19, 0(x0)
    // rom[21] = 32'b000000000010_00000_001_10100_0000011;// lh x20, 2(x0)
    // //rom[x]=32'b imm7  _ rs2 _ rs1 _f3 _ imm5_ op // S-Type
    // rom[22] = 32'b0000000_11111_00010_001_00000_0100011;// sh x31, 0(x2)
    // rom[23] = 32'b0000000_11111_00010_001_00010_0100011;// sh x31, 2(x2)
    // end
    assign data = rom[addr[31:2]];
endmodule
